typedef Int#(8) Input_t;
typedef Int#(16) Output_t;
typedef Int#(32) DTW_Output_t;


typedef 1000   Window_Size;
typedef 8   Input_Size;
typedef 16  Output_Size;
typedef 32  DTW_Output_Size;

typedef 2000  Width;

typedef 4   DivSize;
typedef 4   Module_num;

